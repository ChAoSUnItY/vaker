module vaker

import rand { intn }
import math { pow10 }

const currencies = ['AED', 'AFN', 'ALL', 'AMD', 'ANG', 'AOA', 'ARS', 'AUD', 'AWG', 'AZN', 'BAM',
	'BBD', 'BDT', 'BGN', 'BHD', 'BIF', 'BMD', 'BND', 'BOB', 'BOV', 'BRL', 'BSD', 'BTN', 'BWP',
	'BYN', 'BZD', 'CAD', 'CDF', 'CHE', 'CHF', 'CHW', 'CLF', 'CLP', 'CNY', 'COP', 'COU', 'CRC',
	'CUC', 'CUP', 'CVE', 'CZK', 'DJF', 'DKK', 'DOP', 'DZD', 'EGP', 'ERN', 'ETB', 'EUR', 'FJD',
	'FKP', 'GBP', 'GEL', 'GHS', 'GIP', 'GMD', 'GNF', 'GTQ', 'GYD', 'HKD', 'HNL', 'HRK', 'HTG',
	'HUF', 'IDR', 'ILS', 'INR', 'IQD', 'IRR', 'ISK', 'JMD', 'JOD', 'JPY', 'KES', 'KGS', 'KHR',
	'KMF', 'KPW', 'KRW', 'KWD', 'KYD', 'KZT', 'LAK', 'LBP', 'LKR', 'LRD', 'LSL', 'LYD', 'MAD',
	'MDL', 'MGA', 'MKD', 'MMK', 'MNT', 'MOP', 'MRU', 'MUR', 'MVR', 'MWK', 'MXN', 'MXV', 'MYR',
	'MZN', 'NAD', 'NGN', 'NIO', 'NOK', 'NPR', 'NZD', 'OMR', 'PAB', 'PEN', 'PGK', 'PHP', 'PKR',
	'PLN', 'PYG', 'QAR', 'RON', 'RSD', 'RUB', 'RWF', 'SAR', 'SBD', 'SCR', 'SDG', 'SEK', 'SGD',
	'SHP', 'SLL', 'SOS', 'SRD', 'SSP', 'STN', 'SVC', 'SYP', 'SZL', 'THB', 'TJS', 'TMT', 'TND',
	'TOP', 'TRY', 'TTD', 'TWD', 'TZS', 'UAH', 'UGX', 'USD', 'USN', 'UYI', 'UYU', 'UYW', 'UZS',
	'VES', 'VND', 'VUV', 'WST', 'XAF', 'XAG', 'XAU', 'XBA', 'XBB', 'XBC', 'XBD', 'XCD', 'XDR',
	'XOF', 'XPD', 'XPF', 'XPT', 'XSU', 'XTS', 'XUA', 'XXX', 'YER', 'ZAR', 'ZMW', 'ZWL']

[inline]
pub fn currency(ptr PtrInfo) {
	pointer := &string(ptr.ptr)
	unsafe {
		*pointer = rand_element(vaker.currencies)
	}
}

[inline]
pub fn amount(ptr PtrInfo) {
	amount := precision(rand.f64() * pow10(intn(9) or { 1 }), intn(3) or { 1 } + 1)
	match ptr.sz {
		4 {
			pointer := &f32(ptr.ptr)
			unsafe {
				*pointer = f32(amount)
			}
		}
		8 {
			pointer := &f64(ptr.ptr)
			unsafe {
				*pointer = amount
			}
		}
		else {}
	}
}

[inline]
pub fn amount_with_currency(ptr PtrInfo) {
	amount := precision(rand.f64() * pow10(intn(9) or { 1 }), intn(3) or { 1 } + 1)
	currecy := rand_element(vaker.currencies)
	pointer := &string(ptr.ptr)
	unsafe {
		*pointer = '$amount $currecy'
	}
}

[inline]
fn precision(f f64, pre int) f64 {
	div := pow10(pre)
	return f64(i64(f * div)) / div
}
