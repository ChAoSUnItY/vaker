module vaker

const (
	tld = [
		'com',
		'biz',
		'info',
		'net',
		'org',
		'ru',
		'tw',
		'xyz'
	]
	
)

[inline]
pub fn email(ptr PtrInfo) {
}
